
//
module Input_block(
input clk,
input rst_n,
input button,
input button_sub,
input Mode_sel,
output [8:0]angle_to_show_in,				//传给Show_In_block的角度0-360
output [6:0]angle_to_arith,			//传给Arith_block的角度0-90
output cos_sign_to_output,			//cos符号，传给Show_Out_block
output sin_sign_to_output,				//sin符号，传给Show_Out_block
output c_s_swap_to_output				//cos与sin交换标志，传给Show_Out_block
);



////////////输入角度计数器////////////
//当按钮按下时，开始计数器开始递增//////
reg [25:0]counter_reg;
reg [8:0]temp_angle_to_show;

always@(posedge clk or negedge rst_n) begin
	if(~rst_n) begin 
		temp_angle_to_show <= 0;
		counter_reg <= 0;
	end
	else if(~button) begin								//当按键按下时进行计数
		counter_reg <= counter_reg + 1'b1;			
		if(counter_reg == (26'd5000000)) begin		//计数满5M时，显示数字+1，约为0.1s
			counter_reg <= 0;
			temp_angle_to_show <= temp_angle_to_show + 1'b1;
			if(~Mode_sel && temp_angle_to_show == 360)begin		//不同模式下的最大输入值不同
				temp_angle_to_show <= 9'd0;
			end
			else if(Mode_sel && temp_angle_to_show == 79) begin
				temp_angle_to_show <= 9'd0;
			end
		end
	end
	else if(button_sub) begin
		temp_angle_to_show <= temp_angle_to_show - 1'b1;
	end
end

assign angle_to_show_in = temp_angle_to_show;



reg [8:0]temp_angle_to_arith; 		//临时变量，传递到Arith_block
reg cos_sign; 
reg sin_sign;								//cos 和 sin的正负符号，0表示正，1表示负
reg c_s_swap;								//cos和sin交换标志，0表示不交换，1表示交换

always@(*) begin
		if(temp_angle_to_show >=0 && temp_angle_to_show <= 90) begin
			cos_sign <= 1'b0;											//0-90度，cos为+,sin为+,角度等于显示角度, cos与sin值不交换
			sin_sign <= 1'b0;
			c_s_swap <= 1'b0;
			temp_angle_to_arith <= temp_angle_to_show;
		end
		else if( temp_angle_to_show <= 180) begin
			cos_sign <= 1'b1;											//90-180度，cos为-,sin为+,角度等于显示角度 - 90, cos与sin值交换
			sin_sign <= 1'b0;
			c_s_swap <= 1'b1;
			temp_angle_to_arith <= temp_angle_to_show - 9'd90;
		end

		else if( temp_angle_to_show <= 270) begin
			cos_sign <= 1'b1;											//180-270度，cos为-,sin为-,角度等于显示角度 - 180, cos与sin值不交换
			sin_sign <= 1'b1;
			c_s_swap <= 1'b0;	
			temp_angle_to_arith <= temp_angle_to_show - 9'd180;
		end

		else if( temp_angle_to_show <= 360) begin
			cos_sign <= 1'b0;											//270-360度，cos为+,sin为-,角度等于显示角度 - 270, cos与sin值交换
			sin_sign <= 1'b1;
			c_s_swap <= 1'b1;
			temp_angle_to_arith <= temp_angle_to_show - 9'd270;
		end
end
	
	assign angle_to_arith		= temp_angle_to_arith[6:0]; 
	assign cos_sign_to_output	= cos_sign;
	assign sin_sign_to_output	= sin_sign;
	assign c_s_swap_to_output	= c_s_swap;
/////////////////////////////////////






endmodule


