
module Show_Out_block(



);


endmodule 
